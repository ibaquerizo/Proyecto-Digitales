library ieee;
use ieee.std_logic_1164.all;
USE IEEE.STD_LOGIC_unsigned.ALL;

Entity bit_to_7seg_unidad is
	Port(	w: in std_logic_vector(5 downto 0);
			en: in std_logic;
			Q1: out std_logic_vector(6 downto 0));
end bit_to_7seg_unidad;

Architecture sol of bit_to_7seg_unidad is
Signal F1: std_logic_vector(6 downto 0);

Begin			--gfedcba
	with w select
	F1<=  "1000000"  when "000000"|"001010"|"010100"|"011110"|"101000"|"110010"|"111100", --0 10 20 30 40 50 60
			"1111001"  when "000001"|"001011"|"010101"|"011111"|"101001"|"110011", --1 11 21 31 41 51
			"0100100"  when "000010"|"001100"|"010110"|"100000"|"101010"|"110100", --2 12 22 32 42 52
			"0110000"  when "000011"|"001101"|"010111"|"100001"|"101011"|"110101", --3 13 23 33 43 53
			"0011001"  when "000100"|"001110"|"011000"|"100010"|"101100"|"110110", --4 14 24 34 44 54
			"0010010"  when "000101"|"001111"|"011001"|"100011"|"101101"|"110111", --5 15 25 35 45 55
			"0000010"  when "000110"|"010000"|"011010"|"100100"|"101110"|"111000", --6 16 26 36 46 56
			"1111000"  when "000111"|"010001"|"011011"|"100101"|"101111"|"111001", --7 17 27 37 47 57
			"0000000"  when "001000"|"010010"|"011100"|"100110"|"110000"|"111010", --8 18 28 38 48 58
			"0010000"  when "001001"|"010011"|"011101"|"100111"|"110001"|"111011", --9 19 29 39 49 59
			"1111111"  when others;
	Q1<=not(F1) when en='1' else "0000000"; 
end sol;
